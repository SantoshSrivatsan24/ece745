package i2c_pkg;

    typedef enum bit {WRITE=1'b0, READ=1'b1} i2c_op_t;

endpackage