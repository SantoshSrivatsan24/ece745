import ncsu_pkg::*;

class i2c_transcation extends ncsu_component;


endclass