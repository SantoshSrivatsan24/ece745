import ncsu_pkg::*;

class wb_agent extends ncsu_component;


endclass