class i2cmb_predictor extends ncsu_component #(.T(i2c_transaction));

endclass