class i2c_configuration extends ncsu_configuration;


endclass