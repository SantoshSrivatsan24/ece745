class i2cmb_coverage extends ncsu_component #(.T(i2c_transaction));


endclass