import ncsu_pkg::*;

class wb_monitor extends ncsu_component;

endclass