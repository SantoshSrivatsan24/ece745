class wb_monitor extends ncsu_component #(.T(wb_transaction));

endclass