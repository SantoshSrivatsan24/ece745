import ncsu_pkg::*;

class i2c_agent extends ncsu_component;


endclass