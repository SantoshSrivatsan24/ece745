class wb_agent extends ncsu_component #(.T(wb_transaction));


endclass