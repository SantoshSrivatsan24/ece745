package abc_pkg;

  import ncsu_pkg::*;
  `include "ncsu_macros.svh"

  `include "src/abc_typedefs.svh"
  `include "src/abc_configuration.svh"
  `include "src/abc_transaction_base.svh"
  `include "src/abc_random_transaction.svh"
  `include "src/abc_random_statistics_transaction.svh"
  `include "src/abc_randseq_transaction.svh"
  `include "src/abc_randseq_statistics_transaction.svh"
  `include "src/abc_driver.svh"
  `include "src/abc_monitor.svh"
  `include "src/abc_coverage.svh"
  `include "src/abc_agent.svh"

endpackage
