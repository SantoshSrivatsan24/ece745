class wb_configuration extends ncsu_configuration;


endclass