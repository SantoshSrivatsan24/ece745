class i2cmb_scoreboard extends ncsu_component #(.T(i2c_transaction));

    

endclass