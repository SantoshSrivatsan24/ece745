`define BANNER(t, x) \
	$display ("==========================================================================="); \
	$display ("%s (%t)", x, t); \
	$display ("---------------------------------------------------------------------------");

`define FANCY_BANNER(x) \
	$display ("\n***************************************************************************"); \
	$display ("%s", x); \
	$display ("***************************************************************************\n");