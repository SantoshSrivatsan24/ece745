class i2cmb_generator_fsm_test extends i2cmb_generator_base;

    `ncsu_register_object(i2cmb_generator_fsm_test)

    function new (string name = "", ncsu_component_base parent = null);
        super.new (name, parent);
    endfunction


    virtual task run ();



    endtask

endclass