// `define CSR_ADDR	2'h0
// `define DPR_ADDR 	2'h1
// `define CMDR_ADDR 	2'h2

// `define CMD_START     8'bxxxx_x100
// `define CMD_STOP      8'bxxxx_x101
// `define CMD_READ_ACK  8'bxxxx_x010
// `define CMD_READ_NACK 8'bxxxx_x011
// `define CMD_WRITE     8'bxxxx_x001
// `define CMD_SET_BUS   8'bxxxx_x110
// `define CMD_WAIT      8'bxxxx_x000