class i2cmb_environment extends ncsu_component #(.T(i2c_transaction));

endclass