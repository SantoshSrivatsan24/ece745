import ncsu_pkg::*;

class i2cmb_environment extends ncsu_component;

endclass