import ncsu_pkg::*;

class i2c_monitor extends ncsu_component;


endclass