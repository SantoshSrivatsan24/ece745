package wb_pkg;

    import ncsu_pkg::*;

    `include "src/wb_transaction.svh"
    `include "src/wb_configuration.svh"
    `include "src/wb_agent.svh"
    `include "src/wb_driver.svh"
    `include "src/wb_monitor.svh"

endpackage