class i2cmb_generator extends ncsu_component #(.T(i2c_transaction));

endclass