import ncsu_pkg::*;

class i2c_configuration extends ncsu_component;


endclass