import ncsu_pkg::*;

class i2cmb_test extends ncsu_component;

endclass