import ncsu_pkg::*;

class i2cmb_generator extends ncsu_component;

endclass