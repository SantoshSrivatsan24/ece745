class i2cmb_test extends ncsu_component #(.T(i2c_transaction));

endclass