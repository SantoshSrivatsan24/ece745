import ncsu_pkg::*;

class wb_configuration extends ncsu_component;


endclass