`define BANNER(x) \
	$display ("============================================================"); \
	$display ("%s", x); \
	$display ("------------------------------------------------------------");

`define FANCY_BANNER(x) \
	$display ("\n************************************************************"); \
	$display ("%s", x); \
	$display ("************************************************************\n");

`define SEPARATOR \
    $display ("============================================================");