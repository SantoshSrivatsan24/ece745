import ncsu_pkg::*;

class i2cmb_scoreboard extends ncsu_component;

endclass