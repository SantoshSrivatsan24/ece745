class i2cmb_env_configuration extends ncsu_configuration;

endclass