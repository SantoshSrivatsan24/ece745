import ncsu_pkg::*;

class wb_driver extends ncsu_component;

endclass