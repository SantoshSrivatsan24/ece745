class i2c_agent extends ncsu_component #(.T(i2c_transaction));


endclass