import ncsu_pkg::*;

class i2c_driver extends ncsu_component;


endclass