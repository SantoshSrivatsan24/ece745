package first_project_pkg;

  import ncsu_pkg::*;
  import abc_pkg::*;
  `include "ncsu_macros.svh"

  `include "src/env_configuration.svh"
  `include "src/predictor.svh"
  `include "src/coverage.svh"
  `include "src/scoreboard.svh"
  `include "src/environment.svh"
  `include "src/generator.svh"
  `include "src/test_base.svh"

endpackage
