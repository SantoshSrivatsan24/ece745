import ncsu_pkg::*;

class i2cmb_coverage extends ncsu_component;


endclass