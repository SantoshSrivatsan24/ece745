import ncsu_pkg::*;

class i2cmb_env_configuration extends ncsu_component;

endclass