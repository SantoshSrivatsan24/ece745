import ncsu_pkg::*;

class wb_transaction extends ncsu_component;

endclass