class wb_configuration extends ncsu_configuration;

    function new (string name = "");
        super.new (name);
    endfunction

endclass