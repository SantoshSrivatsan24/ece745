import ncsu_pkg::*;

class i2cmb_predictor extends ncsu_component;

endclass