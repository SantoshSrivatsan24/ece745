class i2c_monitor extends ncsu_component #(.T(i2c_transaction));


endclass