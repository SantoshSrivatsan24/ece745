class i2c_configuration extends ncsu_configuration;

    function new (string name = "");
        super.new(name);
    endfunction
endclass